module registers (RegWrite, WriteRegister, RS, RT, RD, readData1, readData2);
  input RegWrite;
  input [4:0] WriteRegister; //recebe resultado do MUX
  input [4:0] RS; //Read Register 1 parte [25:21] da instrucao
  input [4:0] RT; //Read Register 2 parte [20:16] da instrucao
  input [4:0] RD; //parte [15:11] da instrução
  output [31:0] readData1; //Saida de dados 1
  output [31:0] readData2; //Saida de dados 2

//Banco de registradores
reg [31:0]BancoReg[31:0]; //Armazena dados contidos nos registradores
initial begin
    BancoReg[0] = 32'b00000000000000000000000000000000;
    BancoReg[1] = 32'b00000000000000000000000000000001;
    BancoReg[2] = 32'b00000000000000000000000000000010;
    BancoReg[3] = 32'b00000000000000000000000000000011;
    BancoReg[4] = 32'b00000000000000000000000000000100;
    BancoReg[5] = 32'b00000000000000000000000000000101;
    BancoReg[6] = 32'b00000000000000000000000000000110;
    BancoReg[7] = 32'b00000000000000000000000000000111;
    BancoReg[8] = 32'b00000000000000000000000000001000;
    BancoReg[9] = 32'b00000000000000000000000000001001;
    BancoReg[10] = 32'b00000000000000000000000000001010;
    BancoReg[11] = 32'b00000000000000000000000000001011;
    BancoReg[12] = 32'b00000000000000000000000000001100;
    BancoReg[13] = 32'b00000000000000000000000000001101;
    BancoReg[14] = 32'b00000000000000000000000000001110;
    BancoReg[15] = 32'b00000000000000000000000000001111;
    BancoReg[16] = 32'b00000000000000000000000000010000;
    BancoReg[17] = 32'b00000000000000000000000000010001;
    BancoReg[18] = 32'b00000000000000000000000000010010;
    BancoReg[19] = 32'b00000000000000000000000000010011;
    BancoReg[20] = 32'b00000000000000000000000000010100;
    BancoReg[21] = 32'b00000000000000000000000000010101;
    BancoReg[22] = 32'b00000000000000000000000000010110;
    BancoReg[23] = 32'b00000000000000000000000000010111;
    BancoReg[24] = 32'b00000000000000000000000000011000;
    BancoReg[25] = 32'b00000000000000000000000000011001;
    BancoReg[26] = 32'b00000000000000000000000000011010;
    BancoReg[27] = 32'b00000000000000000000000000011011;
    BancoReg[28] = 32'b00000000000000000000000000011100;
    BancoReg[29] = 32'b00000000000000000000000000011101;
    BancoReg[30] = 32'b00000000000000000000000000011110;
    BancoReg[31] = 32'b00000000000000000000000000011111;
  end
  always @ (WriteRegister) begin
    if(RegWrite == 1'b1) begin
      BancoReg[RD] = WriteRegister;
    end
  end
  assign readData1 = BancoReg[RS];
  assign readData2 = BancoReg[RT];
endmodule